`timescale 1ns/100ps
typedef class Packet;
typedef mailbox #(Packet) pkt_mbox;
